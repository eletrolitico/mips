module cpu(
	input
);

endmodule 