module cpu();

endmodule 