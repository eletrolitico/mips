module instructionmemory(
	input clk,
	input [9:0] addr,
	output reg [31:0] data_out
);

reg [31:0] M[0:1023];
integer k;

initial begin
	M[0] = 32'b0;
	M[1] = 32'b001101_00001_00000_1100_0000_0000_0000; //LW $s0,C000h($s1) ($s0 = $s1 + C000h)
	M[2] = 32'b001101_00010_00001_1100_0000_0000_0001; //LW $s1,C001h($s2) ($s1 = $s2 + C001h)
	M[3] = 32'd0;
	M[4] = 32'd0;
	M[5] = 32'd0;
	M[6] = 32'b001100_00000_00001_00000_01010110010; //MUL $s0,$s1,$s0 ($s0 = $s1*$s0)
	M[7] = 32'b001101_00011_00010_1100_0000_0000_0010; //LW $s2,C002h($s3) ($s2 = $s3 + C002h)
	M[8] = 32'b001101_00100_00011_1100_0000_0000_0011; //LW $s3,C003h($s4) ($s3 = $s4 + C003h)
	M[9] = 32'd0;
	M[10] = 32'd0;
	M[11] = 32'd0;
	M[12] = 32'b001100_00010_00011_00100_01010100000; //ADD $s4,$s2,$s3 ($s4 = $s2+$s3)
	M[13] = 32'd0;
	M[14] = 32'd0;
	M[15] = 32'd0;
	M[16] = 32'b001100_00000_00100_00000_01010100010; //SUB $s0,$s0,$s4 ($s0 = $s0-$s4)
	M[17] = 32'd0;
	M[18] = 32'd0;
	M[19] = 32'd0;
	M[20] = 32'b001110_00101_00000_1100_0011_1111_1111; //SW $s0,C3ffh($s5) (M[$s5 + C3ff] = $s0)
	M[21] = 32'd0;
	M[22] = 32'd0;
	M[23] = 32'd0;
	M[24] = 32'd0; 
	
//PROGRAMA ERRADO
	M[25] = 32'd0;
	M[26] = 32'd0;
	M[27] = 32'd0;
	M[28] = 32'b001101_00111_00110_1100_0000_0000_0000; //LW $s6,C000h($s1) ($s6 = $s7 + C000h)
	M[29] = 32'b001101_01000_00111_1100_0000_0000_0001; //LW $s7,C001h($s8) ($s7 = $s8 + C001h)
	M[30] = 32'b001100_00110_00111_00110_01010110010;   //MUL $s6,$s7,$s6 ($s6 = $s7*$s6)
	M[31] = 32'b001101_01001_01000_1100_0000_0000_0010; //LW $s8,C002h($s9) ($s8 = $s9 + C002h)
	M[32] = 32'b001101_01010_01001_1100_0000_0000_0011; //LW $s9,C003h($s10) ($s9 = $s10 + C003h)
	M[33] = 32'b001100_01000_01001_01010_01010100000;   //ADD $s10,$s8,$s9 ($s10 = $s8+$s9)
	M[34] = 32'b001100_00110_01010_00110_01010100010;   //SUB $s6,$s6,$s10 ($s6 = $s6-$s10)
	M[35] = 32'b001110_01011_00110_1100_0011_1111_1111; //SW $s6,C3ffh($s11) (M[$s11 + C3ff] = $s6)
	for(k = 36; k < 1024; k = k+1) M[k] = 32'b0;
end
	
always @ (posedge clk)
	begin
		data_out <= M[addr];
	end
	
endmodule
